// -----------------------------------------------------------------------------
// ALU Verification — UCF EEE 5703
// Authors: Jonathan Joslin, Patrik Reagan
// Date: 30 November 2024
// -----------------------------------------------------------------------------

class alu_test extends uvm_test;
  `uvm_component_utils(alu_test)
  
  alu_env env;
  alu_test_sequence test_seq;
  
  // Constructo
  function new(string name="alu_test", uvm_component parent);
    super.new(name,parent);
    `uvm_info("TEST_CLASS", "Inside Constructor", UVM_HIGH )
  endfunction: new
  
  // Build Phase
  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    `uvm_info("TEST_CLASS", "Build Phase", UVM_HIGH )

    env = alu_env::type_id::create("env", this);
    
  endfunction: build_phase
  
  // Connect Phase
  function void connect_phase(uvm_phase phase);
    super.connect_phase(phase);
    `uvm_info("TEST_CLASS", "Connect Phase", UVM_HIGH )
    
    // connect monitor with the scoreboard
    

  endfunction: connect_phase

  task run_phase(uvm_phase phase);
    super.run_phase(phase);
    `uvm_info("TEST_CLASS", "Run phase!", UVM_HIGH)
    
    phase.raise_objection(this);
    #10;
    // Start our sequences
    repeat(100) begin
    //test sequence
    test_seq = alu_test_sequence::type_id::create("test_seq");
    test_seq.start(env.agent.sequencer);
    #10;
    end
    phase.drop_objection(this);

    
        
  endtask: run_phase
  
endclass: alu_test